module not1(c, a);
input a;
output c;
assign c=~a;
endmodule